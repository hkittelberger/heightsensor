module rom_8(
    input logic [4:0] col,
    input logic [4:0] row,
    output logic [5:0] data
);

logic [9:0] address;
assign address = {row, col};

    always_comb begin
        case(address)
            10'b0000000000: data = 6'b000000;
            10'b0000000001: data = 6'b000000;
            10'b0000000010: data = 6'b000000;
            10'b0000000011: data = 6'b000000;
            10'b0000000100: data = 6'b000000;
            10'b0000000101: data = 6'b000000;
            10'b0000000110: data = 6'b000000;
            10'b0000000111: data = 6'b000000;
            10'b0000100000: data = 6'b000000;
            10'b0000100001: data = 6'b000000;
            10'b0000100010: data = 6'b000000;
            10'b0000100011: data = 6'b000000;
            10'b0000100100: data = 6'b000000;
            10'b0000100101: data = 6'b000000;
            10'b0000100110: data = 6'b000000;
            10'b0000100111: data = 6'b000000;
            10'b0001000000: data = 6'b000000;
            10'b0001000001: data = 6'b000000;
            10'b0001000110: data = 6'b000000;
            10'b0001000111: data = 6'b000000;
            10'b0001100000: data = 6'b000000;
            10'b0001100001: data = 6'b000000;
            10'b0001100110: data = 6'b000000;
            10'b0001100111: data = 6'b000000;
            10'b0010000000: data = 6'b000000;
            10'b0010000001: data = 6'b000000;
            10'b0010000110: data = 6'b000000;
            10'b0010000111: data = 6'b000000;
            10'b0010100000: data = 6'b000000;
            10'b0010100001: data = 6'b000000;
            10'b0010100110: data = 6'b000000;
            10'b0010100111: data = 6'b000000;
            10'b0011000000: data = 6'b000000;
            10'b0011000001: data = 6'b000000;
            10'b0011000110: data = 6'b000000;
            10'b0011000111: data = 6'b000000;
            10'b0011100000: data = 6'b000000;
            10'b0011100001: data = 6'b000000;
            10'b0011100010: data = 6'b000000;
            10'b0011100011: data = 6'b000000;
            10'b0011100100: data = 6'b000000;
            10'b0011100101: data = 6'b000000;
            10'b0011100110: data = 6'b000000;
            10'b0011100111: data = 6'b000000;
            10'b0100000000: data = 6'b000000;
            10'b0100000001: data = 6'b000000;
            10'b0100000010: data = 6'b000000;
            10'b0100000011: data = 6'b000000;
            10'b0100000100: data = 6'b000000;
            10'b0100000101: data = 6'b000000;
            10'b0100000110: data = 6'b000000;
            10'b0100000111: data = 6'b000000;
            10'b0100100000: data = 6'b000000;
            10'b0100100001: data = 6'b000000;
            10'b0100100110: data = 6'b000000;
            10'b0100100111: data = 6'b000000;
            10'b0101000000: data = 6'b000000;
            10'b0101000001: data = 6'b000000;
            10'b0101000110: data = 6'b000000;
            10'b0101000111: data = 6'b000000;
            10'b0101100000: data = 6'b000000;
            10'b0101100001: data = 6'b000000;
            10'b0101100110: data = 6'b000000;
            10'b0101100111: data = 6'b000000;
            10'b0110000000: data = 6'b000000;
            10'b0110000001: data = 6'b000000;
            10'b0110000110: data = 6'b000000;
            10'b0110000111: data = 6'b000000;
            10'b0110100000: data = 6'b000000;
            10'b0110100001: data = 6'b000000;
            10'b0110100110: data = 6'b000000;
            10'b0110100111: data = 6'b000000;
            10'b0111000000: data = 6'b000000;
            10'b0111000001: data = 6'b000000;
            10'b0111000010: data = 6'b000000;
            10'b0111000011: data = 6'b000000;
            10'b0111000100: data = 6'b000000;
            10'b0111000101: data = 6'b000000;
            10'b0111000110: data = 6'b000000;
            10'b0111000111: data = 6'b000000;
            10'b0111100000: data = 6'b000000;
            10'b0111100001: data = 6'b000000;
            10'b0111100010: data = 6'b000000;
            10'b0111100011: data = 6'b000000;
            10'b0111100100: data = 6'b000000;
            10'b0111100101: data = 6'b000000;
            10'b0111100110: data = 6'b000000;
            10'b0111100111: data = 6'b000000;
            default: data = 6'b111111;
        endcase
    end
endmodule